/**
 * @ Author: German Cano Quiveu, germancq@dte.us.es
 * @ Create Time: 2020-04-14 13:43:32
 * @ Modified by: German Cano Quiveu, germancq
 * @ Modified time: 2022-03-15 15:48:17
 * @ Description:
 */




//////////////////////////////////////////////////////////////////////
///                                                               ////
/// ORPSoC top for Atlys board                                    ////
///                                                               ////
/// Instantiates modules, depending on ORPSoC defines file        ////
///                                                               ////
/// Copyright (C) 2013 Stefan Kristiansson                        ////
///  <stefan.kristiansson@saunalahti.fi                           ////
///                                                               ////
//////////////////////////////////////////////////////////////////////
//// This source file may be used and distributed without         ////
//// restriction provided that this copyright statement is not    ////
//// removed from the file and that any derivative work contains  ////
//// the original copyright notice and the associated disclaimer. ////
////                                                              ////
//// This source file is free software; you can redistribute it   ////
//// and/or modify it under the terms of the GNU Lesser General   ////
//// Public License as published by the Free Software Foundation; ////
//// either version 2.1 of the License, or (at your option) any   ////
//// later version.                                               ////
////                                                              ////
//// This source is distributed in the hope that it will be       ////
//// useful, but WITHOUT ANY WARRANTY; without even the implied   ////
//// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ////
//// PURPOSE.  See the GNU Lesser General Public License for more ////
//// details.                                                     ////
////                                                              ////
//// You should have received a copy of the GNU Lesser General    ////
//// Public License along with this source; if not, download it   ////
//// from http://www.opencores.org/lgpl.shtml                     ////
////                                                              ////
//////////////////////////////////////////////////////////////////////

`include "orpsoc-defines.v"

module orpsoc_top #(
	parameter	rom0_aw = 8,
	parameter	uart0_aw = 3
)(
	input		sys_clk_pad_i,
	input		rst_n_pad_i,



	input next_button,
	input center_button,
	input up_button,
	inout [7:0] gpio0_io,
	output [7:0] leds,
	input [15:0] switch_i,

	//SPI
	output	   sclk,
	output	   mosi,
	input	   miso,
	output 	   cs,
	output SD_RESET,
	output SD_DAT_1,
	output SD_DAT_2,

   // UART
	input		uart0_srx_pad_i,
	output		uart0_stx_pad_o,

	//7seg
	output [6:0] seg,
    output [7:0] AN,
    output DP,

	// DDR2

	output [12:0]	ddr2_addr,
	output [2:0]	ddr2_ba,
	output		ddr2_ras_n,
	output		ddr2_cas_n,
	output		ddr2_we_n,
	output		ddr2_odt,
	output		ddr2_cke,
	output	[1:0]	ddr2_dm,
	inout [15:0]	ddr2_dq,
	inout	[1:0]	ddr2_dqs_p,
	inout	[1:0]	ddr2_dqs_n,
	output      ddr2_cs_n,
	output		ddr2_ck_p,
	output		ddr2_ck_n,


	
	//debug ts
	output inicio_proceso_led,
	output fin_de_proceso_led

);

assign inicio_proceso_led = leds[7];//idle_led from bootloader_module
assign fin_de_proceso_led = leds[6];//finish_led from bootloader_module


parameter	IDCODE_VALUE=32'h14951185;

//SD in SPI_MODE
assign SD_RESET = 1'b0;
assign SD_DAT_1 = 1'b1;
assign SD_DAT_2 = 1'b1;

logic btn_debug;
pulse_button debug_btn_up(
   .clk(wb_clk),
   .reset(1'b0),
   .button(up_button),
   .pulse(btn_debug)
);
////////////////////////////////////////////////////////////////////////
//
// Clock and reset generation module
//
////////////////////////////////////////////////////////////////////////

logic async_rst;
logic wb_clk, wb_rst; //wb_clk generated by ddr
logic dbg_tck;


logic dvi_clk;

logic ddr2_if_clk;
logic ddr2_if_rst;
logic clk100;
logic clk50;
logic clk200;

logic locked_mmcm;
assign ddr2_if_clk = clk200;

dcm_pll_generator clkgen0(
	.global_clk_in(sys_clk_pad_i),
    .rst(~rst_n_pad_i),
    .locked(locked_mmcm),
	.clk200(clk200),
    .clk100(clk100),
    .clk50(clk50)
);



assign clk_bootloader = clk100;


rstgen rstgen0
       (
	// Main clocks in, depending on board
	.sys_clk_pad_i(sys_clk_pad_i),
	// Asynchronous, active low reset in
	.rst_n_pad_i(rst_n_pad_i),
	.locked_mcm(locked_mmcm),

	// Wishbone clock and reset out
	.wb_clk(wb_clk),

	.wb_rst_o(wb_rst),
	.ddr2_if_rst_o(ddr2_if_rst)
);


assign async_rst = ~ rst_n_pad_i;
assign ddr2_clk = ddr2_if_clk;

////////////////////////////////////////////////////////////////////////
//
// Modules interconnections
//
////////////////////////////////////////////////////////////////////////
`include "wb_intercon.vh"





////////////////////////////////////////////////////////////////////////
//
// OR1K CPU
//
////////////////////////////////////////////////////////////////////////

logic	[31:0]	or1k_irq;

logic sig_tick;

logic or1k_rst;

logic boot_cpu_rst;

assign or1k_rst = wb_rst  | boot_cpu_rst  ;

`ifdef OR1200

or1200_top #(.boot_adr(32'hf0000100))
or1200_top0 (
	// Instruction bus, clocks, reset
	.iwb_clk_i			(wb_clk),
	.iwb_rst_i			(wb_rst),
	.iwb_ack_i			(wb_s2m_or1k_i_ack),
	.iwb_err_i			(wb_s2m_or1k_i_err),
	.iwb_rty_i			(wb_s2m_or1k_i_rty),
	.iwb_dat_i			(wb_s2m_or1k_i_dat),

	.iwb_cyc_o			(wb_m2s_or1k_i_cyc),
	.iwb_adr_o			(wb_m2s_or1k_i_adr),
	.iwb_stb_o			(wb_m2s_or1k_i_stb),
	.iwb_we_o			(wb_m2s_or1k_i_we),
	.iwb_sel_o			(wb_m2s_or1k_i_sel),
	.iwb_dat_o			(wb_m2s_or1k_i_dat),
	.iwb_cti_o			(wb_m2s_or1k_i_cti),
	.iwb_bte_o			(wb_m2s_or1k_i_bte),

	// Data bus, clocks, reset
	.dwb_clk_i			(wb_clk),
	.dwb_rst_i			(wb_rst),
	.dwb_ack_i			(wb_s2m_or1k_d_ack),
	.dwb_err_i			(wb_s2m_or1k_d_err),
	.dwb_rty_i			(wb_s2m_or1k_d_rty),
	.dwb_dat_i			(wb_s2m_or1k_d_dat),

	.dwb_cyc_o			(wb_m2s_or1k_d_cyc),
	.dwb_adr_o			(wb_m2s_or1k_d_adr),
	.dwb_stb_o			(wb_m2s_or1k_d_stb),
	.dwb_we_o			(wb_m2s_or1k_d_we),
	.dwb_sel_o			(wb_m2s_or1k_d_sel),
	.dwb_dat_o			(wb_m2s_or1k_d_dat),
	.dwb_cti_o			(wb_m2s_or1k_d_cti),
	.dwb_bte_o			(wb_m2s_or1k_d_bte),

	// Debug interface ports
	.dbg_stall_i			(),
	.dbg_ewt_i			(1'b0),
	.dbg_lss_o			(),
	.dbg_is_o			(),
	.dbg_wp_o			(),
	.dbg_bp_o			(),

	.dbg_adr_i			(),
	.dbg_we_i			(),
	.dbg_stb_i			(),
	.dbg_dat_i			(),
	.dbg_dat_o			(),
	.dbg_ack_o			(),

	.pm_clksd_o			(),
	.pm_dc_gate_o			(),
	.pm_ic_gate_o			(),
	.pm_dmmu_gate_o			(),
	.pm_immu_gate_o			(),
	.pm_tt_gate_o			(),
	.pm_cpu_gate_o			(),
	.pm_wakeup_o			(),
	.pm_lvolt_o			(),

	// Core clocks, resets
	.clk_i				(wb_clk),
	.rst_i				(or1k_rst),

	.clmode_i			(2'b00),

	// Interrupts
	.pic_ints_i			(or1k_irq),
	.sig_tick			(sig_tick),

	.pm_cpustall_i			(1'b0)
);
`endif

`ifdef MOR1KX
mor1kx #(
	.FEATURE_DEBUGUNIT("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.OPTION_ICACHE_BLOCK_WIDTH(5),
	.OPTION_ICACHE_SET_WIDTH(8),
	.OPTION_ICACHE_WAYS(4),
	.OPTION_ICACHE_LIMIT_WIDTH(32),
	.FEATURE_IMMU("ENABLED"),
	.OPTION_IMMU_SET_WIDTH(7),
	.FEATURE_DATACACHE("ENABLED"),
	.OPTION_DCACHE_BLOCK_WIDTH(5),
	.OPTION_DCACHE_SET_WIDTH(8),
	.OPTION_DCACHE_WAYS(4),
	.OPTION_DCACHE_LIMIT_WIDTH(31),
	.FEATURE_DMMU("ENABLED"),
	.OPTION_DMMU_SET_WIDTH(7),
	.OPTION_PIC_TRIGGER("LATCHED_LEVEL"),

	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_RESET_PC(32'h00000100)
) mor1kx0 (
	.iwbm_adr_o(wb_m2s_or1k_i_adr),
	.iwbm_stb_o(wb_m2s_or1k_i_stb),
	.iwbm_cyc_o(wb_m2s_or1k_i_cyc),
	.iwbm_sel_o(wb_m2s_or1k_i_sel),
	.iwbm_we_o (wb_m2s_or1k_i_we),
	.iwbm_cti_o(wb_m2s_or1k_i_cti),
	.iwbm_bte_o(wb_m2s_or1k_i_bte),
	.iwbm_dat_o(wb_m2s_or1k_i_dat),

	.dwbm_adr_o(wb_m2s_or1k_d_adr),
	.dwbm_stb_o(wb_m2s_or1k_d_stb),
	.dwbm_cyc_o(wb_m2s_or1k_d_cyc),
	.dwbm_sel_o(wb_m2s_or1k_d_sel),
	.dwbm_we_o (wb_m2s_or1k_d_we ),
	.dwbm_cti_o(wb_m2s_or1k_d_cti),
	.dwbm_bte_o(wb_m2s_or1k_d_bte),
	.dwbm_dat_o(wb_m2s_or1k_d_dat),

	.clk(wb_clk),
	.rst(or1k_rst),

	.iwbm_err_i(wb_s2m_or1k_i_err),
	.iwbm_ack_i(wb_s2m_or1k_i_ack),
	.iwbm_dat_i(wb_s2m_or1k_i_dat),
	.iwbm_rty_i(wb_s2m_or1k_i_rty),

	.dwbm_err_i(wb_s2m_or1k_d_err),
	.dwbm_ack_i(wb_s2m_or1k_d_ack),
	.dwbm_dat_i(wb_s2m_or1k_d_dat),
	.dwbm_rty_i(wb_s2m_or1k_d_rty),

	.irq_i(or1k_irq),

	.du_addr_i(),
	.du_stb_i(),
	.du_dat_i(),
	.du_we_i(),
	.du_dat_o(),
	.du_ack_o(),
	.du_stall_i(),
	.du_stall_o()
);

`endif

////////////////////////////////////////////////////////////////////////
//
// GENERIC JTAG TAP
//
////////////////////////////////////////////////////////////////////////
/*
wire	dbg_if_select;
wire	dbg_if_tdo;
wire	jtag_tap_tdo;
wire	jtag_tap_shift_dr;
wire	jtag_tap_pause_dr;
wire	jtag_tap_update_dr;
wire	jtag_tap_capture_dr;

tap_top jtag_tap0 (
	.tdo_pad_o			(tdo_pad_o),
	.tms_pad_i			(tms_pad_i),
	.tck_pad_i			(dbg_tck),
	.trst_pad_i			(async_rst),
	.tdi_pad_i			(tdi_pad_i),

	.tdo_padoe_o			(tdo_padoe_o),

	.tdo_o				(jtag_tap_tdo),

	.shift_dr_o			(jtag_tap_shift_dr),
	.pause_dr_o			(jtag_tap_pause_dr),
	.update_dr_o			(jtag_tap_update_dr),
	.capture_dr_o			(jtag_tap_capture_dr),

	.extest_select_o		(),
	.sample_preload_select_o	(),
	.mbist_select_o			(),
	.debug_select_o			(dbg_if_select),


	.bs_chain_tdi_i			(1'b0),
	.mbist_tdi_i			(1'b0),
	.debug_tdi_i			(dbg_if_tdo)
);
*/
////////////////////////////////////////////////////////////////////////
//
// Debug Interface
//
////////////////////////////////////////////////////////////////////////
/*
wire	[31:0]	or1k_dbg_dat_i;
wire	[31:0]	or1k_dbg_adr_i;
wire		or1k_dbg_we_i;
wire		or1k_dbg_stb_i;
wire		or1k_dbg_ack_o;
wire	[31:0]	or1k_dbg_dat_o;

wire		or1k_dbg_stall_i;
wire		or1k_dbg_ewt_i;
wire	[3:0]	or1k_dbg_lss_o;
wire	[1:0]	or1k_dbg_is_o;
wire	[10:0]	or1k_dbg_wp_o;
wire		or1k_dbg_bp_o;
wire		or1k_dbg_rst;

wire		sig_tick;

adbg_top dbg_if0 (
	// OR1K interface
	.cpu0_clk_i	(wb_clk),
	.cpu0_rst_o	(or1k_dbg_rst),
	.cpu0_addr_o	(or1k_dbg_adr_i),
	.cpu0_data_o	(or1k_dbg_dat_i),
	.cpu0_stb_o	(or1k_dbg_stb_i),
	.cpu0_we_o	(or1k_dbg_we_i),
	.cpu0_data_i	(or1k_dbg_dat_o),
	.cpu0_ack_i	(or1k_dbg_ack_o),
	.cpu0_stall_o	(or1k_dbg_stall_i),
	.cpu0_bp_i	(or1k_dbg_bp_o),

	// TAP interface
	.tck_i		(dbg_tck),
	.tdi_i		(jtag_tap_tdo),
	.tdo_o		(dbg_if_tdo),
	.rst_i		(wb_rst),
	.capture_dr_i	(jtag_tap_capture_dr),
	.shift_dr_i	(jtag_tap_shift_dr),
	.pause_dr_i	(jtag_tap_pause_dr),
	.update_dr_i	(jtag_tap_update_dr),
	.debug_select_i	(dbg_if_select),

	// Wishbone debug master
	.wb_rst_i	(wb_rst),
	.wb_clk_i	(wb_clk),
	.wb_dat_i	(wb_s2m_decoy_dat),
	.wb_ack_i	(wb_s2m_decoy_ack),
	.wb_err_i	(wb_s2m_decoy_err),

	.wb_adr_o	(wb_m2s_decoy_adr),
	.wb_dat_o	(wb_m2s_decoy_dat),
	.wb_cyc_o	(wb_m2s_decoy_cyc),
	.wb_stb_o	(wb_m2s_decoy_stb),
	.wb_sel_o	(wb_m2s_decoy_sel),
	.wb_we_o	(wb_m2s_decoy_we),
	.wb_cti_o	(wb_m2s_decoy_cti),
	.wb_bte_o	(wb_m2s_decoy_bte)
);
*/

////////////////////////////////////////////////////////////////////////
//
// ROM
//
////////////////////////////////////////////////////////////////////////

assign	wb_s2m_rom0_err = 1'b0;
assign	wb_s2m_rom0_rty = 1'b0;

`ifdef BOOTROM
rom #(.addr_width(rom0_aw))
rom0 (
	.wb_clk		(wb_clk),
	.wb_rst		(wb_rst),
	.wb_adr_i	(wb_m2s_rom0_adr[(rom0_aw + 2) - 1 : 2]),
	.wb_cyc_i	(wb_m2s_rom0_cyc),
	.wb_stb_i	(wb_m2s_rom0_stb),
	.wb_cti_i	(wb_m2s_rom0_cti),
	.wb_bte_i	(wb_m2s_rom0_bte),
	.wb_dat_o	(wb_s2m_rom0_dat),
	.wb_ack_o	(wb_s2m_rom0_ack)
);
`else
assign	wb_s2m_rom0_dat_o = 0;
assign	wb_s2m_rom0_ack_o = 0;
`endif


////////////////////////////////////////////////////////////////////////
//
// BOOTLOADER MODULE
//
////////////////////////////////////////////////////////////////////////


logic ram0_mux;




logic ram0_ack;
logic ram0_rst;
logic ram0_we;
logic ram0_cyc;
logic ram0_stb;
logic ram0_cti;
logic [3:0] ram0_sel;
logic [31:0] ram0_data;
logic [31:0] ram0_addr;
logic [31:0] bootloader_debug_data;

/*
bootloaderModule boot0(
	.wb_clk	(wb_clk),
	.wb_rst (center_button),
	.start (1'b1),
	.cpu_rst (boot_cpu_rst),

	.wb_ack_i(wb_s2m_bootloader_ack),
	.wb_we_o(wb_m2s_bootloader_we),
	.wb_cyc_o(wb_m2s_bootloader_cyc),
	.wb_stb_o(wb_m2s_bootloader_stb),
	.wb_sel_o(wb_m2s_bootloader_sel),
	.wb_dat_o(wb_m2s_bootloader_dat),
	.wb_adr_o(wb_m2s_bootloader_adr),

	.mosi(mosi),
	.miso(miso),
	.sclk(sclk),
	.cs(cs),

	.sclk_speed(switch_i[11:8]),
	.cmd_18(switch_i[15]),

	.finish_signal (fin_de_proceso_led),
    .debug_leds (leds[3:0]),
	.debug_sw(switch_i[1:0]),
	.debug_data (bootloader_debug_data)

);
*/

logic [63:0] exec_timer;

wb_raw_boot #(
	.WB_DATA(32),
	.SDSPI_WB_ADDR(32'h92000000),
	.RAM_WB_ADDR(0)
)
boot0(
	.wb_clk(wb_clk),
	.wb_rst(wb_rst),
	.wb_ack_i(wb_s2m_bootloader_ack),
	.wb_err_i(wb_s2m_bootloader_err),
	.wb_dat_i(wb_s2m_bootloader_dat),
	.wb_rty_i(wb_s2m_bootloader_rty),
	.wb_dat_o(wb_m2s_bootloader_dat),
	.wb_cyc_o(wb_m2s_bootloader_cyc),
	.wb_stb_o(wb_m2s_bootloader_stb),
	.wb_sel_o(wb_m2s_bootloader_sel),
	.wb_we_o (wb_m2s_bootloader_we),
	.wb_cti_o(wb_m2s_bootloader_cti),
	.wb_bte_o(wb_m2s_bootloader_bte),
	.wb_adr_o(wb_m2s_bootloader_adr),


	.start(1'b1),
	.cpu_rst(boot_cpu_rst),
	.start_block(32'h0),
	.total_blocks((1<<14)), //8MB/512 2^(23-9) - 1
	.sclk_speed(4'h1),
	.debug(bootloader_debug_data[15:0]),
	.exec_timer(exec_timer),
	.btn_dbg(btn_debug)
);


////////////////////////////////////////////////////////////////////////
//
// ELUKS MODULE
//
////////////////////////////////////////////////////////////////////////

wb_sdspi #(
	.CLK_FQ_KHZ(100000)
) wb_sdspi_inst(
	.wb_clk(wb_clk),
	.wb_rst(wb_rst),
	.wb_adr_i(wb_m2s_sdspi0_adr),
	.wb_dat_i(wb_m2s_sdspi0_dat),
	.wb_we_i (wb_m2s_sdspi0_we),
	.wb_cyc_i(wb_m2s_sdspi0_cyc),
	.wb_stb_i(wb_m2s_sdspi0_stb),
	.wb_sel_i(wb_m2s_sdspi0_sel),
	.wb_cti_i(wb_m2s_sdspi0_cti),
	.wb_bte_i(wb_m2s_sdspi0_bte),
	.wb_ack_o(wb_s2m_sdspi0_ack),
	.wb_err_o(wb_s2m_sdspi0_err),
	.wb_rty_o(wb_s2m_sdspi0_rty),
	.wb_dat_o(wb_s2m_sdspi0_dat),
	.sclk(sclk),
	.cs(cs),
	.mosi(mosi),
	.miso(miso),
    .debug(bootloader_debug_data[31:16])
);


////////////////////////////////////////////////////////////////////////
//
// DDR2 SDRAM Memory Controller
//
////////////////////////////////////////////////////////////////////////

//clock period 200Mhz
//controller operates at 200Mhz/4 = 50Mhz
xilinx_ddr2 xilinx_ddr2_0 (
	.wbm0_adr_i	(wb_m2s_ddr2_bus_adr),
	.wbm0_bte_i	(wb_m2s_ddr2_bus_bte),
	.wbm0_cti_i	(wb_m2s_ddr2_bus_cti),
	.wbm0_cyc_i	(wb_m2s_ddr2_bus_cyc),
	.wbm0_dat_i	(wb_m2s_ddr2_bus_dat),
	.wbm0_sel_i	(wb_m2s_ddr2_bus_sel),
	.wbm0_stb_i	(wb_m2s_ddr2_bus_stb),
	.wbm0_we_i	(wb_m2s_ddr2_bus_we),
	.wbm0_ack_o	(wb_s2m_ddr2_bus_ack),
	.wbm0_err_o	(wb_s2m_ddr2_bus_err),
	.wbm0_rty_o	(wb_s2m_ddr2_bus_rty),
	.wbm0_dat_o	(wb_s2m_ddr2_bus_dat),

	.wb_clk		(wb_clk),
	.wb_rst		(wb_rst),

	.ddr2_addr		(ddr2_addr[12:0]),
	.ddr2_ba	(ddr2_ba),
	.ddr2_ras_n	(ddr2_ras_n),
	.ddr2_cas_n	(ddr2_cas_n),
	.ddr2_we_n	(ddr2_we_n),
	.ddr2_odt	(ddr2_odt),
	.ddr2_cke	(ddr2_cke),
	.ddr2_dm	(ddr2_dm[0]),
	.ddr2_udm	(ddr2_dm[1]),
	.ddr2_ck_p	(ddr2_ck_p),
	.ddr2_ck_n	(ddr2_ck_n),
	.ddr2_dq	(ddr2_dq),
	.ddr2_dqs_p	(ddr2_dqs_p[0]),
	.ddr2_dqs_n	(ddr2_dqs_n[0]),
	.ddr2_cs_n  (ddr2_cs_n),
	.ddr2_udqs_p	(ddr2_dqs_p[1]),
	.ddr2_udqs_n	(ddr2_dqs_n[1]),
	.ddr2_if_clk	(ddr2_if_clk),
	.ddr2_if_rst	(ddr2_if_rst)
);

////////////////////////////////////////////////////////////////////////
//
// GPIO 0
//
////////////////////////////////////////////////////////////////////////

logic [7:0]	gpio0_in;
logic [7:0]	gpio0_out;
logic [7:0]	gpio0_dir;

// Tristate logic for IO
// 0 = input, 1 = output
genvar                    i;
generate
	for (i = 0; i < 8; i = i+1) begin: gpio0_tris
		assign gpio0_io[i] = gpio0_dir[i] ? gpio0_out[i] : 1'bz;
		assign gpio0_in[i] = gpio0_dir[i] ? gpio0_out[i] : gpio0_io[i];
	end
endgenerate

gpio gpio0 (
	// GPIO bus
	.gpio_i		(gpio0_in),
	.gpio_o		(gpio0_out),
	.gpio_dir_o	(gpio0_dir),
	// Wishbone slave interface
	.wb_adr_i	(wb_m2s_gpio0_adr[0]),
	.wb_dat_i	(wb_m2s_gpio0_dat),
	.wb_we_i	(wb_m2s_gpio0_we),
	.wb_cyc_i	(wb_m2s_gpio0_cyc),
	.wb_stb_i	(wb_m2s_gpio0_stb),
	.wb_cti_i	(wb_m2s_gpio0_cti),
	.wb_bte_i	(wb_m2s_gpio0_bte),
	.wb_dat_o	(wb_s2m_gpio0_dat),
	.wb_ack_o	(wb_s2m_gpio0_ack),
	.wb_err_o	(wb_s2m_gpio0_err),
	.wb_rty_o	(wb_s2m_gpio0_rty),

	.wb_clk		(wb_clk),
	.wb_rst		(wb_rst)
);



////////////////////////////////////////////////////////////////////////
//
// UART0
//
////////////////////////////////////////////////////////////////////////

logic	uart0_irq;

uart_top uart16550_0 (
	// Wishbone slave interface
	.wb_clk_i	(clk50),
	.wb_rst_i	(wb_rst),
	.wb_adr_i	(wb_m2s_uart0_adr[uart0_aw-1:0]),
	.wb_dat_i	(wb_m2s_uart0_dat),
	.wb_we_i	(wb_m2s_uart0_we),
	.wb_stb_i	(wb_m2s_uart0_stb),
	.wb_cyc_i	(wb_m2s_uart0_cyc),
	.wb_sel_i	(4'b0), // Not used in 8-bit mode
	.wb_dat_o	(wb_s2m_uart0_dat),
	.wb_ack_o	(wb_s2m_uart0_ack),

	// Outputs
	.int_o		(uart0_irq),
	.stx_pad_o	(uart0_stx_pad_o),
	.rts_pad_o	(),
	.dtr_pad_o	(),

	// Inputs
	.srx_pad_i	(uart0_srx_pad_i),
	.cts_pad_i	(1'b0),
	.dsr_pad_i	(1'b0),
	.ri_pad_i	(1'b0),
	.dcd_pad_i	(1'b0)
);

////////////////////////////////////////////////////////////////////////
//
// 7 seg
//
////////////////////////////////////////////////////////////////////////
logic [31:0] debug_7_seg;
display #(.N(32),.CLK_HZ(100000000)) seg7(
    .clk(wb_clk),
	.rst(wb_rst),
	.din(debug_7_seg),
	.seg(seg),
	.an(AN)
);
//assign debug_7_seg = switch_i[15] ? wb_m2s_or1k_i_adr : wb_s2m_or1k_i_dat;//bootloader_debug_data;
assign debug_7_seg = switch_i[15]==1 ? exec_timer[63:32] : exec_timer[31:0];//{bootloader_debug_data[15:0],4'b0,1'b0,wb_s2m_sdspi0_ack,wb_m2s_sdspi0_cyc,wb_m2s_sdspi0_stb,1'b0,wb_s2m_ddr2_bus_ack,wb_m2s_ddr2_bus_cyc,wb_m2s_ddr2_bus_stb};

////////////////////////////////////////////////////////////////////////
//
// Interrupt assignment
//
////////////////////////////////////////////////////////////////////////

assign or1k_irq[0] = 0; // Non-maskable inside OR1K
assign or1k_irq[1] = 0; // Non-maskable inside OR1K
assign or1k_irq[2] = uart0_irq;
assign or1k_irq[3] = 0;
assign or1k_irq[4] = 0;
assign or1k_irq[5] = 0;
assign or1k_irq[6] = 0;
assign or1k_irq[7] = 0;
assign or1k_irq[8] = 0;
assign or1k_irq[9] = 0;
assign or1k_irq[10] = 0;
assign or1k_irq[11] = 0;
assign or1k_irq[12] = 0;
assign or1k_irq[13] = 0;
assign or1k_irq[14] = 0;
assign or1k_irq[15] = 0;
assign or1k_irq[16] = 0;
assign or1k_irq[17] = 0;
assign or1k_irq[18] = 0;
assign or1k_irq[19] = 0;
assign or1k_irq[20] = 0;
assign or1k_irq[21] = 0;
assign or1k_irq[22] = 0;
assign or1k_irq[23] = 0;
assign or1k_irq[24] = 0;
assign or1k_irq[25] = 0;
assign or1k_irq[26] = 0;
assign or1k_irq[27] = 0;
assign or1k_irq[28] = 0;
assign or1k_irq[29] = 0;
assign or1k_irq[30] = 0;
assign or1k_irq[31] = 0;

endmodule : orpsoc_top // orpsoc_top
